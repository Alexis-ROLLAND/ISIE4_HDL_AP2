module chronometre(ClkIn, DigitH, DigitL);

input ClkIn;

output[0:6] DigitH, DigitL;





endmodule 
